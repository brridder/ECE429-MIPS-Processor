// Memory implementation

module mem{
	   clock,
	   address,
	   data,
	   wren,
	   q
};
   