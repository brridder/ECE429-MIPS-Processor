//
// ALU function definitions
//

`ifndef _alu_func_vh_
`define _alu_func_vh_

`define ADD  6'b100000
`define ADDU 6'b100001
`define SUB  6'b100010
`define SUBU 6'b100011
`define SLT  6'b101010
`define SLTU 6'b101011
`define SLL  6'b000000
`define SRL  6'b000010
`define SRA  6'b000011
`define AND  6'b100100
`define OR   6'b100101
`define XOR  6'b100110
`define NOR  6'b100111

`endif