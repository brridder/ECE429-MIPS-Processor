//
// Control register constant definitions
//

`ifndef _control_vh_
`define _control_vh_

`define CONTROL_REG_SIZE 4

`define REG_WE 0
`define I_TYPE 1
`define R_TYPE 2
`define J_TYPE 3

`endif 
