//
// Control register constant definitions
//

`ifndef _control_vh_
`define _control_vh_

`define CONTROL_REG_SIZE 2
`define REG_WE 0
`define R_TYPE 1

`endif 
