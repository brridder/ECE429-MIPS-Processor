//
// Control register constant definitions
//

`ifndef _control_vh_
`define _control_vh_

`define CONTROL_REG_SIZE 1
`define REG_WE 0

`endif 
